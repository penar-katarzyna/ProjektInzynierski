LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY LCD_display IS
PORT(
	CLK		: IN STD_LOGIC
	
);
END LCD_display;

ARCHITECTURE behavior of LCD_display IS

BEGIN

PROCESS 
BEGIN
WAIT UNTIL(CLK'EVENT) AND (CLK = '1');
END PROCESS;

END behavior;