library IEEE;
use IEEE.STD_LOGIC_1164.all;

package chars is

type LCD_CHARS is array (1 to 2, 1 to 16) of std_logic_vector(7 downto 0);

end chars; 

package body chars is


end chars; 
